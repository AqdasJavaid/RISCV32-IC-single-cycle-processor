
/* ALU Arithmetic and Logic Operations
----------------------------------------------------------------------
|ALU_Sel |   ALU Operation
----------------------------------------------------------------------
| 0  |   ALU_Out = A + B;
----------------------------------------------------------------------
| 1  |   ALU_Out = A - B;
----------------------------------------------------------------------
| 2  |   ALU_Out = A ^ B;
----------------------------------------------------------------------
| 3  |   ALU_Out = A | B;
----------------------------------------------------------------------
| 4  |   ALU_Out = A & B;
----------------------------------------------------------------------
| 5  |   ALU_Out = A << B;
----------------------------------------------------------------------
| 6  |   ALU_Out = A >> B;
----------------------------------------------------------------------
| 7  |   ALU_Out = A >>> B;
----------------------------------------------------------------------
| 8  |   ALU_Out = A < B; //slt
----------------------------------------------------------------------
| 9  |   ALU_Out = unsigned A < unsigned B; //sltu
----------------------------------------------------------------------
| 10  |   ALU_Out = rs2 << 12; //lui
----------------------------------------------------------------------
| 11  |   ALU_Out = pc + (rs2 << 12); //auipc
----------------------------------------------------------------------*/
//

module alu #(parameter width = 32)(
    input wire signed [width-1:0]rs1,
    input wire signed [width-1:0]rs2,
	input wire [3:0]alu_sel,

    output reg [width-1:0]rd

);

always@(*)
	begin
		case(alu_sel)
			4'd0: rd = rs1 + rs2;  //add
			4'd1: rd = rs1 - rs2;  //sub
			4'd2: rd = rs1 ^ rs2;   //xor
			4'd3: rd = rs1 | rs2;   //or
			4'd4: rd = rs1 & rs2;   //and
			4'd5: rd = rs1 << rs2;  //sll
			4'd6: rd = rs1 >> rs2;  //srl
			4'd7: rd = rs1 >>> rs2; //sra
			4'd8: rd = rs1<rs2;     //slt
			4'd9: rd = ($unsigned (rs1)<$unsigned (rs2)); //sltu
			4'd10: rd = rs2;//{rs2[19:0],{12{1'b0}}};   		  //lui
			//4'd11: rd = rs1 + {rs2[19:0],{12{1'b0}}};     //auipc

		default: rd=32'd0;
		endcase
	end

endmodule



